configuration mc8051_datamux_rtl_cfg of mc8051_datamux is

  for rtl
    
  end for;

end mc8051_datamux_rtl_cfg;
