configuration mc8051_clockdiv_rtl_cfg of mc8051_clockdiv is

  for rtl
    
  end for;

end mc8051_clockdiv_rtl_cfg;
