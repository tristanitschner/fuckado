configuration mc8051_chipsel_rtl_cfg of mc8051_chipsel is

  for rtl
    
  end for;

end mc8051_chipsel_rtl_cfg;
